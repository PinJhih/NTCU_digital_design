module Top(
    input [3:0]sw,
    input [3:0]dip_pin,
    output [5:0]led
);
    bin_adder adder(num1,num2, sum);

endmodule
